<?xml version="1.0" encoding="UTF-8" standalone="no"?>
<!-- Created with Inkscape (http://www.inkscape.org/) -->

<svg
   width="48.000004mm"
   height="297mm"
   viewBox="0 0 48.000004 297"
   version="1.1"
   id="svg1"
   xmlns="http://www.w3.org/2000/svg"
   xmlns:svg="http://www.w3.org/2000/svg">
  <defs
     id="defs1" />
  <g
     id="layer1">
    <path
       style="fill:none;stroke:#000000;stroke-width:1.265;stroke-linecap:round;stroke-dasharray:none;stroke-opacity:1"
       d="m 2.3195691,11.218688 c 0,0 7.0328,16.247593 3.34759,37.474859 -3.31832,19.113908 16.9829309,37.413816 12.5223809,59.002573 -3.51033,16.98972 -16.9081309,15.43952 -14.5736609,48.57381 1.1158,15.83705 -1.1536,13.49326 1.92604,59.31816 3.70956,55.19805 4.09556,69.88759 4.16043,70.73094"
       id="path1" />
  </g>
</svg>
